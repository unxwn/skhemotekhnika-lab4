library verilog;
use verilog.vl_types.all;
entity Ex_Polishchuk is
    port(
        x3              : in     vl_logic;
        x2              : in     vl_logic;
        x1              : in     vl_logic;
        f1              : out    vl_logic;
        f2              : out    vl_logic
    );
end Ex_Polishchuk;
